module obstacle #(
    parameter CIDXW=3,
    parameter CORDW=10
    ) (
        input CLK;
        input RESET;
        input line,
        input [3:0] state,
        input [9:0] hc,
        input [9:0] vc,
    );

endmodule